module WriteToMIF;
    reg [15:0] new_data; // New data to be written
    reg [15:0] memory [0:255]; // 16-bit memory with 256 entries

endmodule