

module ArduinoAdd_p1(input logic [19:0] arduinoAdd, output logic [19:0] arduinoAddO);


	assign arduinoAddO = arduinoAdd + 1;


endmodule