
module probe_pc (
	probe);	

	input	[31:0]	probe;
endmodule
